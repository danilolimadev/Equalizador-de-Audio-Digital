module converter_Q5_8 ( 
    input [7:0] gain_in,
    output reg [12:0] gain_out
);
    always @* begin 
        case (gain_in)
            6'b000001:
                gain_out = 13'b00000_00010000; // 1/16
            6'b000010:
                gain_out = 13'b00000_00010001; // 1/15
            6'b000011:
                gain_out = 13'b00000_00010010; // 1/14
            6'b000100:
                gain_out = 13'b00000_00010100; // 1/13
            6'b000101:
                gain_out = 13'b00000_00010101; // 1/12
            6'b000110:
                gain_out = 13'b00000_00010111; // 1/11
            6'b000111:
                gain_out = 13'b00000_00011010; // 1/10
            6'b001000:
                gain_out = 13'b00000_00011100; // 1/9
            6'b001001:
                gain_out = 13'b00000_00100000; // 1/8
            6'b001010:
                gain_out = 13'b00000_00100101; // 1/7
            6'b001011:
                gain_out = 13'b00000_00101011; // 1/6
            6'b001100:
                gain_out = 13'b00000_00110011; // 1/5
            6'b001101:
                gain_out = 13'b00000_01000000; // 1/4
            6'b001110:
                gain_out = 13'b00000_01010101; // 1/3
            6'b001111:
                gain_out = 13'b00000_10000000; // 1/2
            6'b010000:
                gain_out = 13'b00001_00000000; // 1
            6'b010001:
                gain_out = 13'b00001_00000000; // 0 -> 1
            6'b010010:
                gain_out = 13'b00001_00000000; // 1
            6'b010011:
                gain_out = 13'b00010_00000000; // 2
            6'b010100:
                gain_out = 13'b00011_00000000; // 3
            6'b010101:
                gain_out = 13'b00100_00000000; // 4
            6'b010110:
                gain_out = 13'b00101_00000000; // 5
            6'b010111:
                gain_out = 13'b00110_00000000; // 6
            6'b011000:
                gain_out = 13'b00111_00000000; // 7
            6'b011001:
                gain_out = 13'b01000_00000000; // 8
            6'b011010:
                gain_out = 13'b01001_00000000; // 9
            6'b011011:
                gain_out = 13'b01010_00000000; // 10
            6'b011100:
                gain_out = 13'b01011_00000000; // 11
            6'b011101:
                gain_out = 13'b01100_00000000; // 12
            6'b011110:
                gain_out = 13'b01101_00000000; // 13
            6'b011111:
                gain_out = 13'b01110_00000000; // 14
            6'b100000:
                gain_out = 13'b01111_00000000; // 15
            6'b100001:
                gain_out = 13'b10000_00000000; // 16
            default:
                gain_out = 13'b00000_00000000;
        endcase
    end
endmodule
